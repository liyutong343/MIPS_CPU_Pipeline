// 待修改！�??
`timescale 1ns / 1ps
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	initial begin
	   Instruction <= 32'h0;
	end
	
	always @(*)
		case (Address[9:2])
        8'd0: Instruction <= 32'h24050000;
        8'd1: Instruction <= 32'h24070200;
        8'd2: Instruction <= 32'h00002020;
        8'd3: Instruction <= 32'h00054021;
        8'd4: Instruction <= 32'h8d090000;
        8'd5: Instruction <= 32'h11200003;
        8'd6: Instruction <= 32'h20840001;
        8'd7: Instruction <= 32'h21080004;
        8'd8: Instruction <= 32'h08100004;
        8'd9: Instruction <= 32'h00003020;
        8'd10: Instruction <= 32'h00074021;
        8'd11: Instruction <= 32'h8d090000;
        8'd12: Instruction <= 32'h11200003;
        8'd13: Instruction <= 32'h20c60001;
        8'd14: Instruction <= 32'h21080004;
        8'd15: Instruction <= 32'h0810000b;
        8'd16: Instruction <= 32'h00042080;
        8'd17: Instruction <= 32'h00063080;
        8'd18: Instruction <= 32'h0c100036;
        8'd19: Instruction <= 32'h3044000f;
        8'd20: Instruction <= 32'h0c10004c;
        8'd21: Instruction <= 32'h00034021;
        8'd22: Instruction <= 32'h35080e00;
        8'd23: Instruction <= 32'h304400f0;
        8'd24: Instruction <= 32'h00042102;
        8'd25: Instruction <= 32'h0c10004c;
        8'd26: Instruction <= 32'h00034821;
        8'd27: Instruction <= 32'h35290d00;
        8'd28: Instruction <= 32'h30440f00;
        8'd29: Instruction <= 32'h00042202;
        8'd30: Instruction <= 32'h0c10004c;
        8'd31: Instruction <= 32'h00035021;
        8'd32: Instruction <= 32'h354a0b00;
        8'd33: Instruction <= 32'h3044f000;
        8'd34: Instruction <= 32'h00042302;
        8'd35: Instruction <= 32'h0c10004c;
        8'd36: Instruction <= 32'h00035821;
        8'd37: Instruction <= 32'h356b0300;
        8'd38: Instruction <= 32'h3c014000;
        8'd39: Instruction <= 32'h34240010;
        8'd40: Instruction <= 32'hac880000;
        8'd41: Instruction <= 32'h0c100031;
        8'd42: Instruction <= 32'hac890000;
        8'd43: Instruction <= 32'h0c100031;
        8'd44: Instruction <= 32'hac8a0000;
        8'd45: Instruction <= 32'h0c100031;
        8'd46: Instruction <= 32'hac8b0000;
        8'd47: Instruction <= 32'h0c100031;
        8'd48: Instruction <= 32'h08100028;
        8'd49: Instruction <= 32'h24100000;
        8'd50: Instruction <= 32'h241130d4;
        8'd51: Instruction <= 32'h22100001;
        8'd52: Instruction <= 32'h1611fffe;
        8'd53: Instruction <= 32'h03e00008;
        8'd54: Instruction <= 32'h24080000;
        8'd55: Instruction <= 32'h24090000;
        8'd56: Instruction <= 32'h24020000;
        8'd57: Instruction <= 32'h00865022;
        8'd58: Instruction <= 32'h0148082a;
        8'd59: Instruction <= 32'h1420000f;
        8'd60: Instruction <= 32'h24090000;
        8'd61: Instruction <= 32'h0126502a;
        8'd62: Instruction <= 32'h11400008;
        8'd63: Instruction <= 32'h01095020;
        8'd64: Instruction <= 32'h01455020;
        8'd65: Instruction <= 32'h8d4a0000;
        8'd66: Instruction <= 32'h00e95820;
        8'd67: Instruction <= 32'h8d6b0000;
        8'd68: Instruction <= 32'h154b0002;
        8'd69: Instruction <= 32'h21290004;
        8'd70: Instruction <= 32'h0810003d;
        8'd71: Instruction <= 32'h15260001;
        8'd72: Instruction <= 32'h20420001;
        8'd73: Instruction <= 32'h21080004;
        8'd74: Instruction <= 32'h08100039;
        8'd75: Instruction <= 32'h03e00008;
        8'd76: Instruction <= 32'h20010000;
        8'd77: Instruction <= 32'h10240020;
        8'd78: Instruction <= 32'h20010001;
        8'd79: Instruction <= 32'h10240020;
        8'd80: Instruction <= 32'h20010002;
        8'd81: Instruction <= 32'h10240020;
        8'd82: Instruction <= 32'h20010003;
        8'd83: Instruction <= 32'h10240020;
        8'd84: Instruction <= 32'h20010004;
        8'd85: Instruction <= 32'h10240020;
        8'd86: Instruction <= 32'h20010005;
        8'd87: Instruction <= 32'h10240020;
        8'd88: Instruction <= 32'h20010006;
        8'd89: Instruction <= 32'h10240020;
        8'd90: Instruction <= 32'h20010007;
        8'd91: Instruction <= 32'h10240020;
        8'd92: Instruction <= 32'h20010008;
        8'd93: Instruction <= 32'h10240020;
        8'd94: Instruction <= 32'h20010009;
        8'd95: Instruction <= 32'h10240020;
        8'd96: Instruction <= 32'h2001000a;
        8'd97: Instruction <= 32'h10240020;
        8'd98: Instruction <= 32'h2001000b;
        8'd99: Instruction <= 32'h10240020;
        8'd100: Instruction <= 32'h2001000c;
        8'd101: Instruction <= 32'h10240020;
        8'd102: Instruction <= 32'h2001000d;
        8'd103: Instruction <= 32'h10240020;
        8'd104: Instruction <= 32'h2001000e;
        8'd105: Instruction <= 32'h10240020;
        8'd106: Instruction <= 32'h2001000f;
        8'd107: Instruction <= 32'h10240020;
        8'd108: Instruction <= 32'h240300ff;
        8'd109: Instruction <= 32'h0810008e;
        8'd110: Instruction <= 32'h240300c0;
        8'd111: Instruction <= 32'h0810008e;
        8'd112: Instruction <= 32'h240300f9;
        8'd113: Instruction <= 32'h0810008e;
        8'd114: Instruction <= 32'h240300a4;
        8'd115: Instruction <= 32'h0810008e;
        8'd116: Instruction <= 32'h240300b0;
        8'd117: Instruction <= 32'h0810008e;
        8'd118: Instruction <= 32'h24030099;
        8'd119: Instruction <= 32'h0810008e;
        8'd120: Instruction <= 32'h24030092;
        8'd121: Instruction <= 32'h0810008e;
        8'd122: Instruction <= 32'h24030082;
        8'd123: Instruction <= 32'h0810008e;
        8'd124: Instruction <= 32'h240300f8;
        8'd125: Instruction <= 32'h0810008e;
        8'd126: Instruction <= 32'h24030080;
        8'd127: Instruction <= 32'h0810008e;
        8'd128: Instruction <= 32'h24030090;
        8'd129: Instruction <= 32'h0810008e;
        8'd130: Instruction <= 32'h24030088;
        8'd131: Instruction <= 32'h0810008e;
        8'd132: Instruction <= 32'h24030083;
        8'd133: Instruction <= 32'h0810008e;
        8'd134: Instruction <= 32'h240300c6;
        8'd135: Instruction <= 32'h0810008e;
        8'd136: Instruction <= 32'h240300a1;
        8'd137: Instruction <= 32'h0810008e;
        8'd138: Instruction <= 32'h24030084;
        8'd139: Instruction <= 32'h0810008e;
        8'd140: Instruction <= 32'h2403008e;
        8'd141: Instruction <= 32'h0810008e;
        8'd142: Instruction <= 32'h03e00008;


			
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
